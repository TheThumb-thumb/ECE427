import le_types::*;
import params::*;
module oht_tb;

logic clk, rst;

initial clk= 1'b0;
always #1ns clk= ~clk;
initial rst= 1'b0;

    logic adc_in, deque;
    logic perm_fail, valid;
    logic [7:0] calibration_arr_n, calibration_arr_p;
    // logic clk_div;
    logic [1023:0] input_val;
    logic [9:0] counter;

    always_ff @(posedge clk) begin
        if (rst) begin
            adc_in <= '0;
            input_val <= 1024'b0000000000000000000000000000000111111111111111111111111111111100000000000000000000000000000001111111111111111111111111111111000000000000000000000111111111111111111111000000000000000000000111111111111111111111111111111100000000000000000000000000000001111111111111111111111111111111000000000000000000000111111111111111111111111111111100000000000000000000011111111111111111111111111111110000000000000000000000000000000111111111111111111111000000000000000000000111111111111111111111111111111100000000000000000000000000000001111111111111111111111111111111000000000000000000000000000000011111111111111111111111111111110000000000000000000001111111111111111111111111111111000000000000000000000111111111111111111111111111111100000000000000000000000000000001111111111111111111110000000000000000000001111111111111111111111111111111000000000000000000000111111111111111111111111111111100000000000000000000011111111111111111111111111111110000000000000000000001111111111111111111111111111111000000000000000000000111111111111111111111000000;
            counter <= '0;
        end else begin
            adc_in <= input_val[counter];
            counter <= counter + 1;
        end
    end

    OHT dut (
        .adc_in(adc_in),
        .clk(clk),
        .rst(rst),
        .debug_mode(1'b0),
        .spi_reg_lsb('0),
        .full(1'b0),
        .perm_fail(perm_fail),
        .valid(valid),
        // calibration output
        .calibration_arr_n(calibration_arr_n),
        .calibration_arr_p(calibration_arr_p)
    );

    initial begin
		$fsdbDumpfile("oht_dump.fsdb");
		$fsdbDumpvars(0, "+all");
		rst = 1'b1;
        #10ns
		rst = 1'b0;
		#100000ns
		$finish();
	end


endmodule