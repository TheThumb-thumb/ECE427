import uvm_pkg::*;

module top_tb;
    

endmodule
