import le_types::*;
import params::*;
module oht_top_tb;

logic clk, rst;

initial clk = 1'b0;
always #1ns clk = ~clk;
initial rst = 1'b0;

    logic [es_sources-1:0] ES_in; // 0-31 latch 32-63 jitter
    logic deque;                  // tells us aes is reading? Does that matter?
    logic debug_mode;
    logic [15:0] spi_reg_lsb;

    logic [cond_width-1:0] cond_out;
    logic full;
    logic empty;
    logic [latch_sources-1:0][calib_bits-1:0] arr_n;
    logic [latch_sources-1:0][calib_bits-1:0] arr_p;
    logic [jitter_sources-1:0] j_disable_arr;
    logic [es_sources-1:0] rd_good_arr;

    logic [1023:0] test_vec [0:100];

    assign test_vec[0] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign test_vec[1] = 1024'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign test_vec[2] = 1024'b0000000000000000000000000000000000000000000000000000000100000010000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000001000000000000000010000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000;
    assign test_vec[3] = 1024'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000001010000100000000000000000000000001000000000000100000000000000000000000000000000000000100000000101000100000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000010000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000000000000000001000000000000000100000000000000000000000000000000000100000000000000000000000000101000000000000100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000;
    assign test_vec[4] = 1024'b0000000000000000000001000000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000001000000100000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001000000000000000000001000000000100000000001000000000000000000000000100000000000000000000000000000000000001000001000100000000000001000000000010000000000000000000000000000000000000000100000000001110000000000000000000000000001000000000000000000000000001000001000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000010000100000000000000001000000000000000000000000100000000000000000000000000000010000000000000000000001000000000000000000000001000000000000000000000000000000000010000000000000000000000000001000000000000000001100000000000000000000000000000000000000000;
    assign test_vec[5] = 1024'b0000000000000000000000000000000000000000000000001000000000000000001000000000000000000000100000000000010010000000000000000000000000010000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000010000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000100000000010000000000001000000000000000000000000001000000100000100000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000001000000000000000000000100000001000000001000000000000000000000000000000000101001000010010010000000000000000000000000000011100000000000000000000100000000100000000001001100000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000100000000000000000000000010000000000000000000000001000000010000000000000000100000000000000000000000000000001000000000000000000000100000000000000000000000100000000;
    assign test_vec[6] = 1024'b0000000011000000000010000000000000000000000001000000000000000000000001100000000000000000000011000000000000000000000000000000000000100000001000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000100000000000000000000001000000000000000000000000000000000000010000000001000000000000100000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000010000000000000000000100000000000000000000000001000100000010000000010000000000000000100100000011110000000000001100000000000000000000100000000000000000000000010000001000000000000000000000000001000000001000000000001000000001000100001000000010010000010000010000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000000000000000001000000000000100001000000000100000000000000000000000000000000000000000010100000000000000000000100000000000000100000000010000;
    assign test_vec[7] = 1024'b0000000000000100001000000000000010000001000000000000001010110000000000010000000000000000000000000000000011000000000101100000000000000000000000000000000000000000000000000000000001000000000001000000010000000000000000001000000000000000110100010001001100000000001010000000000000000001010000000001001000010000000000000000000000000000000000000000000000010000000000000000000000100000000000000000001100010000000000000000000000000101000000000010000000100000000000000000000000000010000001100000000010000000000000000000000100000000000000000000000110000000000000000000000000010000001000000000000000100000000000000000000000000000000000000000001000000000000000000000000000000100100000000000001000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000000000001000000000000000000000000000000000100000000000000000100000000000000000000000000000010000000000000000000000100000000000000000000000000000000000100001000000000100010000000000000100010000000001;
    assign test_vec[8] = 1024'b0000000000000010000000000000000000000000000010100000001000000010000000001000000000000010000010000000000000001000101000001000000000000010001000000000000000010000100001001100001010000001010000000000001000000000000000000000000100000100000000001000000000000000001000000000100100100000000000000000001000000000000000001000101100000000000000000010000000000000000001000000000000101000000000010000000000000000100010000000000000000000000000000000000000000000000001000000000000000000000000000001000000000100000000000000000100000000000000100000000000000000000000000000000000000000000001000000000000000000000000000010000000000000000001000110000000000000000000000010000000000000000000000000001000100000000000001000000000000000000000000010000000010000000000001001000000000000000000000000000000010000000000000000011000000000000010000000000000000000001011000000000000000001000000000000000110001000000000000000000011000000000000000000000000000000100000000000000000000000001000000000000000000000001000100010000001000000000000000001000000000000;
    assign test_vec[9] = 1024'b0010000000000000000000000000000000000001000000000100001000000000000000010000000000000100000000000100000000000000010010000000100000000100010001010000100000000000000000000000001000000000000100001000000000000001000000010010000010000100100100000000000000000000000010000000000100000000000000000000100000000000001000000000100000000010000000000010000010000000000000000000000000000000000000000000000000000001100000000000000000000000000000010000101000000000010000000000000100000100000000001000100000001000000000001000100000000000000000000000000000000100100000000000000000000011000000000001000000000000000000000000010000100000000000000000110001000000100000001000000000000000000000000000001000010000000000100000010000000000000001000000000000000001100010000100001000010000000000000001000000000000001000000000001001000000000000000000000100100100000001100000000000000000000100000000000000001000010000000000010000000000000000000000000001000000000000000000000011110000000000001000000000000000001000100000000000010000000000001000000000000000;
    assign test_vec[10] = 1024'b0000000000000100000000000010000000000000000000010001000000000000000000000000010000011010100000000000000000000000000000001000000000000000100000000000000000001000000000000110000000000010000000000000000100000001000000100000001000000000000000000000000010010001000000000000001001000000001100000000000001000000000010000010000000001000001000000010000100010100000000100000011000100000010010001000000001000000000000000011000000000000010000000001000000000000000000000000000000000101000000000000010000000000000000000000000000000100000000000000000100000001000000000100100001000000000000000000000001001000000000000100000001100000001000100010000000010111001000000000000010000100000000100000000000001000000000000001000000000000000100000000000000100000000000000000000000000000000001000000000000000010000000000000110000000000000000000010100000000100000000000000000001000000000001010000000000000010000000000000000000000000000000000000000000000000000100001000010001000000000100000000000000100100010010000000001000001000000000001000010101000000;
    assign test_vec[11] = 1024'b0000000000000000000001010000000000000000100010100000000100000001000000000101000000000000000010000000000001000000000000110000001000100100000000010000000011000100010000000000100000000010000001001000000000000000010100000000000000001000001000000000000000000010000000000000100000010010000000000000000000000000000000000000000000000000010010000000000000001100001000000001000000000001000001000010000000010000010000000000000000010000001000000000110000000000011000000000000000000000000010000001000000000000100010000000000010000000000000000000000000000000000001100000000000001001000100000010000000000010000011000001000000000000000000000000000001001000000100100000101000100000100000000000000000000100000000000000000000000001001000010000010000000100000000000100000000100001000010000000000000000101001000000000000100001000010000000010000000000100000000000000000001000000110100001000001000000100000100000100001010000100000000000000000000000000000000011000000000000100000000000000000000000000000110001000000000011000000000000010000000000000;
    assign test_vec[12] = 1024'b0000000000000000000010000000000000100000000000000010100000000000000000000000100010000100000000001000001000000100000000001000000000000000000000000000000110100000100000000000000000100010000000000000010000001000001001000000000101000000000001000000000000001000001000000000010000000010000000000010000000000000000000000000000010010000000100000000000000000010000000000100001000001001000000000000000000000100001000000000010000000001001100000000000001001000000000000000001000010010000000100001010000000001000000010011000000100000000000100000001000011001000000001000001001000000000000000000100000000001000000000000000100001000001000000000000011000000000000100001101000000100000010000000001000000000101010010000000000101110000000000000000000101000001000001000000000000000000000001000000000100000010001000000000100000000000010010001000000100000100000000000000001000000101000000000100100000000001000000010000001000111000000001000000000101000000100000000000000000000000000000000001000001000010000000000000001000010000000100000000000000100;
    assign test_vec[13] = 1024'b0000100000010000100000100000000000010000001101000010001000000000100100000000000001100000100000000000001001000000000010000000000000000000011000000001000000000000010000000000000000100000000000000000000000000000000000001000000000000010000000001000010000100000000010010000110010000000100001000000000000000000001000110000000010000101000100001001100000000010000010000000000100000000100000001000000000000000110000000000000000100000000000000000000000010000000100000000000100000001000000101100000000000000000001000000000000000000000000101000010010000000000001000100000000000100000001000010010000100010000000000000100000110000100110100000000000010000000000000000000000100000000000000001000000000000100000001010000000000000000000000000000000001000000000000100000001001011000000000000100000000001000000000011000001001001100001000000000100000000000010001000100000010000100000000100000000110001100011000000011001000000000000010000000000000000000001000100000000000000000000000000100000101000000000000000100101100110001010010000000000000100;
    assign test_vec[14] = 1024'b0000010100000000001000000000010000000001000100000000000100010000001000000000010000000000001000000000001000000000001000010001001000000000000110000010000010000001000000000000000010000000000001001000000000100000101010000000010000001110000000000101100100000000100010001001000001010010000100000000000000000000010000000100000010000100000001000000000000000000000001100000001001000100000000100010000010000000000100010000000100000100000000001001001000000001000000000000000101000000001100001001000000000000000010010010000000000000000000010000000000000011001000000000000100100000000000000000000100000000000000000100000000000000010110000100000000000000100000010000000101000000010001010000010000000110000000000001100000001000000000001000000000000100000000110000000000010000100000000000000000000000000000000000000000001000100000011000000000010000000000000000000000010000001000000000110010000010000000001010100100100001000100000010000000100000000011000010000000000011000100100100000000001000001010001000100001001000000000010000000000010100;
    assign test_vec[15] = 1024'b0000000000001001001000010000010000001001010010001000000000000100000000000000000000100000001000100000000001000001000000000000001000000000000000000000001000000001011000001000000000000000000000000000000000000000100000000000011001000001001000101010011000010000010000000000100010000000100100011000010010000000000000010010001000000000100100000010000010010000000000000000000000001001000000100000000000100000000101000000100000000000001010010010000101000000100001000000000010001100001101000000000000011000000011100110000000000010010000000001010000000000000000000000110001101010000000100000000001010001000100000000000010100000000000000001010001000000001100001001000000000000000000101001000000010010000000000110000000000000000000000100100000001000000000000000000001000000100000000001000000000001000000101010000000000010000010000000000000110100100000000010000000000000011001010000000000000100000000000000000001000000000010000000001000001000100010110000100000001100001000000000001100000101000000010000000000000100100000000100000100000000;
    assign test_vec[16] = 1024'b0000100010000000100000000000000000010000000000000000000100000000000000000000100000100010100000101110000100010000010000000101100000100010000010000000010110000010000001001100100001000000000000110000001100000100000001001101001100000000000000010010000001000010000010000000101000011000011000010100110000011000000001001110000100001000001000000010000010000000010000000010100100000000000100000000000000100000000000100100000000000000000100000010000000001101000001010110000000000000000000000000100000001000100100000001100010000100000110000000000010010100010000011000001010001000000000100000000110100000010000000010000001010100000000000000000000010010000010000001100000001000100100000000000000000000000000000000000000000000000000000000100100000000010100000000000010000110000011000000000000000000000000001000100000000001100010000000000000000000000000000000000000000110000010000001000000001011000001001000100000010000010100000000001010000000000010000000010100010001000100100000000100000000000000000000000010100000000000000000010000100010;
    assign test_vec[17] = 1024'b0000000000010010110011010000000000100000010010001011000010110010011010000000101011000000100010000000001100000001101100100000011000000000001000000000000001011001000000000000000000001001010000100101000000100000001101000110000001001010000001000100001100001000000000000000000001000000000100000000000000000100010100000000100010000010000000000000100100000000000000000000000001000000000000000000000001000010011000000100100010000010000000000000001000010000001100001001010000000001000000000000001001000110011001000010010000000000000000100000000000000101000010000000010000001000000000000000000101000100001000101001100000001001000001000011000100000000000001010000000100001100000101000000100000100000000111101000000000100010010000010000001000000000001100000100000101000000000000000000000001001000000000000000000000000000000010001000100000100100000100000000001001000000100000000000000000000000000000010010001000100000000000000000100100000100010000000000000000110001000000000110001001000000010000001000100001110000000000000010000000100000;
    assign test_vec[18] = 1024'b0101000000100000000001010100010000000000000000000000000001000000000100011000000100001000001000010000010010000000000100000000001100000001100000101000000010001010000001100000000010010100000000010000001000000010000001000100010000000010000000011000000000000000111100010000011100111000001100100000100000110000000001000000000000000001010111000000000000000000001001100000000000100000000000000010101100100000000000010000100001001000110100000000000100000010100101100000000000001011100000000000000000000000001010010001000000010000100101100100000000100000000001000010100000000000010000000000000011001100110011111100000001000000000001000000001100000010000000000000001100000011000010000000011000100011010000000000010010001000000100000001000000000100000010000000000000001000000011010000000100000001100000000100001110000000001010100000010001001000010000010000000100000010000000100010000000010000101011000101000000000000100000100010101000000000010000000000000000000100001000000001010001010000000000000000001000000000000000000000000000100000;
    assign test_vec[19] = 1024'b0000000000010001010100000100000000001000100000100000000100100000000000000100000001010110000000101000000011001000100000001101001000000001000000011000000000000000100000000101110010000000000101010000001000000100101000000000010011010000000000010000001000000000001010001100000001110001001010000000000000000000000000100000000000000110000010000000000000010010000010001000000000000000100000000101000001000010000100000000000000000010001010110000111000010100000000010001000000100001000001010001000010001000001000000001000010100000000110000111000000000110000001011010010000100001100000110001010001001001001110010000000000000000010011001001100010000000100001000001000010010000000000100010000000001000010100000100000001000000100000001110101010000001000000000100000000001001000000110000101100000000010000000110000001010100100001010100000011100000000000000000000000101000100000000000000100001000100001011000000100000000001000000000000000100000010001000100100101000000000000100000000000000000010000000000010000000000000000100011000010000100;
    assign test_vec[20] = 1024'b0000000010000001001001000100000000000011000000000000000000001000001001000001000101001000100000000010010100011000000001000000000000111000000000000110100101000000000000001000101000000000000000000000000000000000101100000011010010000000001000001010000000000000000100101011001010010000000000000000000000000011101110000010000100000010000000101000000000000001000010001000000000000011000000000010010000001000100000001001001010001001000000010011100001000000000000000100000000000010001110010000000010010011100000000111100000000110101010100101100001110000000101000000000101001000010000000000100010000000000100000000100100000000101000110100000000101000100000001000000000000010000110101100100000010110010000000001001011000100011000010000110000010101100010000101000101001000000000000000100010001000001000011000000000000100000000001000000000100000001110000000101000100000000101000000000000000000000010000000000100001000100000000010010100100000000000000000000110010000010101000000001000110010010000010000000100000010100110000000011000001000;
    assign test_vec[21] = 1024'b0000001000000000000000001000000000000011100000000000000101001000101001000000010000010000001000000000000000100000000001010100000100000100001000000000100100100100000000101010100001010100000000001000000100010000001000000100001010101110001010000000010010100000100000010000000010000001000000000000010001111000100100000000000010000000000010100001001000000010000000101110000001000000000000000000000010100010001000110000001000000000000000000000000000110000000000010100101011000000000000101101000000100010001011000000001010000000111000100010010001001010101000000011000001000010000000101000000000000001100001011010110000100001001101000010001000000100010101000000000110000011001000000100000100001000010011000000000100100110010101000000000100000011001010001010110000000000000000010001000010000000010000101011000100000000000100110100000000110110101000001111000000100000100010001000000010010000000000000000000000000110000010000001000100000100100000001011000000010101000000000000000100000110010111100001000000000010000000000100000011000001;
    assign test_vec[22] = 1024'b0001000001000100000011000110001000000000100000010100000010100010100000000100000100000000000000000100110000001000010000000001000000000010111010000000000001000001100110101010001000010011001000000000010101000000011000000010000011100000010000000100000000000000000000000000000000000000010000010000000001001000001000011000000000101000011001001011000001000000000001000100000000101010000100100101110000011100000100100000000101100110001000110000100010010000011000010000001000110000000010100000010000010001101110010010000010111000001000100001101001000110001001000000010000100110001000000000111000000000100000000010000011001000101101000000111000000000001100000000010000000010001010000000010001001101000100110000000000000001000100000000000000100000001000011000110000001000010000000001000000000110011000010000011000000000101010000000010000100101110001001000000000100001010000001000000000000000010000011101000000000011001100100000000111000000100010000000000000000010000100001000101000010110001001000000000011000000000001000000100001011000;
    assign test_vec[23] = 1024'b0000100000000010010000000011000110100001101100100000011001000000100000000000000010000001000000000000010000000110010000001000000010000000000000000001010001000010001000001001001000001010100101011010100000000000101000000110010000001010010100000110100010001010110000001001001000000000110010001000100001111000000000010100010010000000100001100001001001100000100010000001001010000101001001001000011011010010000000010000010000010001000001001100001001001000100000100100100100000000111110000001001000001000000010111000100000000100001100010010010001100010011000000000000010100001000000011100010001000001000000100000000000001000000101001000001000001100100000000010110100000100000011000000000000010100000100000000110110000000000000001001101000001010000001000100001100010110000000010010010000000000100000000001001100010001100100101110000010000000000000000000100000011000000111100000000111000000010000100000000000100001000010100000100000111000010000010000000010000000000000001110000000000000100100000001110000101000000100000100000010001000;
    assign test_vec[24] = 1024'b1000100101000001101001000100000011000000000000100001001110010000111100000000000000000010000010000000001000000110010100100100010011100100000110010000000001100100001000000100101111000001100110000000000011010000001110000000111010000100000100000000000001000000100001000010110000000000010010101010100000101101000100101000000000001000001101000000001000010010010000010001000101100000000000000001100100000000000000100011001001010011001000000000000001010000000000000011100100000010011000000000000000000000000010001000000000100000000110001000010000000000010000100100110001000000001011010000010100010000000000001000000001010000000000000000000111100001001000011000100000001000001010101100001110000000010101010010010001001000001000100010100010001000000000100000001010001001100000000100010110100100000000000010101000010101010000110000000100010011100100000000001100101001000100000100110000000100010000001000010010001000000010000100011100110000000111011000001000001000100100000001000001000000000000010000010000001001000011010011011000100010;
    assign test_vec[25] = 1024'b0000000000000000000010010000001010000000101000100100000000000100100000011000110001000000000000100110001000000000000110010001110000001000010011000100000000000010000000000000100000011001011011110000000101100000101000000111011000000010010101001000010001000000001100111001000100000001010000000000010100001000000001001000010001000000010000000001000000010001101000111001100100000010111010000000001010000100100010010000110010000001100010010001011000001000110000000010110000010000011000011100110100001010000100110000000010000000101000000000100011100110000111000000000101000010111010100011100000000010000000010000001000001100010010000000001100000000000111011100000000000010000000000000001000011110000000000001001101000000001000000010001011100000001001010000000100000001000000000010001111000001000000010000111010010110001000010000001001000000100000010010001010100000001010100100010001100000001000010101110101000000100000000000100101100000000001101101000110110100001100100000000110011000001010000100000000000000010000001101010000000010;
    assign test_vec[26] = 1024'b0000001000110000000011001000100000000000010100001001100101010000001001001011101000010110000000000101100000000101010010011000110001000010001000011000100000010000110011100010000001010010001000000011001001000001000001101010000100000110011000111000011000011010011000010101110010001010000101100010000000000001100001110000000111111001010000010101100010011000000000010001001000000101000000011100000000000000000000111010000110000011000000110001001000011101000110110010000101000000010000000100011100000001101000100100101000000000001000001001000111000000000100010101000000000000101000000110001100000000011000100000000000000010111100101100101010000000100101000100001010100000000001000010101000000000000010010000100000000000000100010000000100000001000000000000000010011100000001000000000010100010101000110101001011000001010011110000000000110100000011001000000100101000001010000000000001000010100000000000000000010100010000001000010010001001000010001110001001001000000000010000000001000001110001000010011000001000000100101000000000010000;
    assign test_vec[27] = 1024'b1001010011010000001001001000010111101000110011101010001000100000000000001100010000000100000110001000000000100000010001000111000010010001000001100110000000010000000000000100100100010000010100000000100010001100100000000000011010000000101000010011001000011100000001001001010000101000000000001110000010010110010000010011100100000110100000000001001100000100001010000001100000001000100000111100000000000010000001001010001110001000101100000100110100010000000100110000101010010000100000110001011101000001000110001000011001010001010100000010000010000110000000000000101101000000100010010100000000111010000001010000100010001010000001000010000000010001010000001101010111000010000100011011101000000100110010000010000101000111010001110000001000000000000000001001010001110100111000000100010000010111000010000001000000100100100110000001100001010100100001000000000010001100010000010000000010001000000100000001111100001010000000110000000010110000000000000000011001000000011000000110110110000011011000000001000100000000010000010010000101010000;
    assign test_vec[28] = 1024'b0100001110000001110000110000011110000110010011000001000100101000101000000110010000010111001000011100000101011011100011110000100100110000000000000001001110000100000110001100100001001000100101001000110100100100010000010000001000010000000000000000011000000110110001000110010011001000000000000010011000110000000101001010011000100010110110010011001110000000000000000110000001000000001010000101000000000001010100001000000100000001100100000011001101000000001000000100010001110100010111001000100001010000001000100011000010001000110000000001000011000000010000111110010000000001010000000110001100101001000001010000111101000101010001001101000001100000000001101100000001010000001000001010000100000000010010000000001100100000100001001000000010100110000011110100011010010010000101000100000100001011001101000100100000000000001000100000001001100100000010000100111100100101100000000000000100001101001000101010000100000000101000001000000100100000101001000001100011110000000000000001000010011100000000000000001011001000000011100000001100000000;
    assign test_vec[29] = 1024'b0111101000100010010001011001000011010100000100001010010011001100000000100000001100000000101100001110100011001001010001000000100000011000111011010000011000101010010000100000010011001011000010011001010100010000100000000000000011110000000010000010101000011010001000010100001001000000001000000000110100010010001000100001010010011011001000000000000000101100100100111000000001001001000000100001100001000011010010001000001110010100011011011110010000101011000001000010110100111000000001001100001000100011000000100110000101110100000010001011000000100110000010000110100100010000001011100000000000000000010100000010100001010100001000001100011000011110000001001000101011110000000000100100000010000000000000000000001010100000000010100001100110011010100000001000001000000000000000101001010100000111010000000010000001101000000010001111010000110011010000000001000011111000000000010010100011000001100010000000000000000110001000000011000000000001000110000100001000000010000110001100110100000000110000110010010100010100000001110011000000101011;
    assign test_vec[30] = 1024'b0111100000010001010100000000000101110000011001100000001100010100100101100010000000000101100011010110010100001111000000110010000001010000010110001010010110100100000101010000100101001001100110011100100000010001000100101100000111101000100000000100001000100000001111010011001001000010000100001000000000000001000000000110101000011100000001000100000010000000010110111000000010010011000000000010000011010011000101000001001001100011000001001000001000111001001011010000000000000000100100101001000000000001000011000100000001001010000100101100010110001010101010100110000100001000100101101000001011010010011010010011100001010100000011010001010000000001010000000000001000000100100000011000110000101011100100011100010101001010010000000001100111000010000000001001011000000010001001001000101000100101110011000011000101100010000000001010000000100010000010000010100001000000001010000011011001010000000000101110000001100010111111000001000000000000010110101000000000010001011000000010111111000110010010000001000001000001000010010000000111000000;
    assign test_vec[31] = 1024'b0100101100000011000001000111010000101000000111000010001010100110011111101100000100000000101001110001000000110000001100100010001001000000010010011000000001011100000001010100100000011011000001000000000010001000110100111010001001011000011000100100001000110010011101101100000011000010000110110010100100010000100101101101000010111100000000000100100000110000001001000001000010011011010000010100000010110010000110000110100000001000000000010000001001000000000001111010010000001100010100110100100010101000001100001000000010110000000000110000000100011110000001000111100011100110010110110001000000000111110000000010010001001001010000000000000000100011000100110010100111001100110001000100000100000001000001101001000000011110000000000111010110001000000000001000011100000000000000100010110100001000000010100111001001100101000000000100000000101011010101010100101001000000010000110010000010100000010011000011000110000000100110100010010000010010101000110000001001101010000010100011000110010010001111000000010010010110000000000010000100110010;
    assign test_vec[32] = 1024'b0100001000100100011000000001010000000000000001010010010000111000000000001100000010111001001010101000011001101010001010100010011100000010000001111110000001001000000000001000100110011000001110000000100000001001010001010100111000000110000011010101000001100000110101101011001000000101001100011010000111010000110100100101001100001000010000000101010000001111010000001000100001000010001001110101001100100001000100000010101011000001000001110010110000100010011100100000000010110000001100000001000000000010111001000101100000101101010010100001001110000101001101010010100100010010001110001010000101000010010111111000001001101000010100010000000011000010001011001000000010000000001001001001000001000001000000010010010001000010010000111001010101100110000100011000101010100100001000000000100010100110011001000110000001010010100000010111000001010001001000001001100001100000010000011000011110001011001010000100100100010000010000000100010111011110100001000111110000011010011101000011000100001100001100100000010000000100010000010011000001000010;
    assign test_vec[33] = 1024'b0100100000100011100001110000001100110000010001011000101110100110011000101100010000000000011000000101010010000100000100000011000001110101001000110100100000011000100010100111100010000000011000000110011010101001010000010110101000001001000011000111010001101000011001100111000011001010011101000110001101010011100100001100000010110010011010100000011001010010010010000110001100010000000001001001000101000010011001000010000000100100001100000101000101000101001100001011000110010000000010001100100001100001100010100000000011001000110000010110000010101000101100111111100011000000111000000011000000101000100001111000000000111011000000110100000100010111010000011000011001100000000000010010000100110100000000100100000001000000100000101000000010000100001100000000010001000010000000010111011001000000010100000110100000000011100011000011000001000100000000000001001010101010000100010011001000010111000010000110000101000001001001000100010011111100100100010001110011100010000000001110110001010101100011100010000001000001001110100011010001111110;
    assign test_vec[34] = 1024'b0001101001001110011100100100000001000110101100011000000000010001000110011100001110000000000000101000101000001100000100000100000001001101100001000000000001110001110001000111100000000100010000000010000000100010010011000001110100100000100110001101100010011011001001100000010001000001100100101000100011101011000011100111010000011000101100000011010000000101010000010011010001010010100100100000100101101010100000010101111000110101010100000010100000110011100000001100010011011101000000110000000000100000101000100000000000011001000000000111010001010100101001001001010010000101000000010101000011000010001000010000101100000001101000000001010000000000000001011010000011110000011000011100100010000000010010010110100100010011010101010110000001001110000010100011010001010100010010111111010110001110010101010110100001111011100001011001000001110010111111010100101010100110001000000100010000101010110001110010000100001011101000010000100111000010000000000000110000100100010011011111001110001100000001000110000001100001011100000000011000110000;
    assign test_vec[35] = 1024'b0000110000101000111001101100001000000000010100100110011100010101011111010001001010100100101010000010000101011000100100000110110010001111000100110010101010100110100111111010000011001000101101010111000011011100011010100100011000010000001010101001100011000110101000010000100010000000010001110000110010000001100110100000100000000000001101010001001000001000100000010001001000100100100110110011100101010010000000100000110100111010110000000111001000110000110100001011110010000000010100000010110110110011001000111001010100000010000101000010110000101111010001011001110010010001000010010011001100001000011000010000111100000001010001000010010010100100111110001000011000010000000100100000000100010011100000000000101001001001100001101010001100000011010001011001010100001000000000000000010000100000111011000001100001000010001000111100010010100000001100111001100100100010000010001110000010111001000101011001000010010001010000101010101000100000001000010100110001111101000001110000010001010000010000000000010011110000001001100100010100111100;
    assign test_vec[36] = 1024'b1100001000011010100001101100101011000101000101000000100000111010011001011000101100001101001000001001001010011000101000000000011000001000010011010100100000100111000001011100110110010010100001101011011010010000000001000011000001100000011011001000000100011001010001011100100000100010001000000110010111101000011001000000110001000001110101111010100010010111001101100111101001010101100100110010100011100000011011000000100001110011001000001000000010000110000001101110110000010000000001101101110000100000110101000010010000000100000110100110101100000100000010111011100001000001010101001001101111000100010100100101111010000001001100010111100110000010000111011000010101000010001001000010001010110010111001010000100100000000000001000001010100100000101110110010111100110011000111110000000000011001000000000000100010111110010000000000000010010101101010100001101001010100101111111001010100110100000101111000000110010000100100010100000000000000000000000111100000001001100001110000001001001100010100000001101001010000010100101000001101100100;
    assign test_vec[37] = 1024'b0010010100100110100100000101000101001110000000000001000110110010010000000010000010010111011010000011000110111011001000000100010000011100010001100001000001000000000001110011000101110101000011100100011010100001110100000011001110010000000101000100001000100101000011100110001000110000010010001000101000111001000000011001000000000000101110010100010001011111011111110110100000100000111100110111100001000001000001100000000010100001010001110000011011000010110110001110001101100000000000111000011001100001000100011011010001001010000100000010101100000010010001010000010000000011001100101110010010110100001000010101000111001000010101111101011110100110110100001010000110100111011010011111110010110001100101000100010101011000011100010101110110001100010111000001111000100100111000011100011010001010010000000001110000100000010101000000111010101100000010010010000110001000000100010000000000000001000000001101001110010001000111100110100001010010110000011000100110001000000101101000110001000010101001001101101110010000001101001101100011000011;
    assign test_vec[38] = 1024'b1000010110010000100011010000000111100100100001110000010001011010000000001010010010100010000100011000011111100000010010111110111000011100010010001010000000000000100010100100110100001111011110000000101000110100110000101011010001110001001110000000101101101000000011011111100011100100001000011101001000000000100111001101001010000101111011000010001001001010000110000001111101001001001000000101000000001100010011111101000001010000011110000111100010010011000000101101001000000110101000110000010100100100000100111000100100000110100100100011010101011100111100110011100000000001101001100111101111000110000110000000000010111111001000000100010100000001001000011011100110000101111010101001100011000010001011000111000000000101010001000111011000000001110000111010000100000011000110000000000010110110001001001010100010010100101010111000011101111010010010001000010101111001111001010001100000110100001010110011010000000000011001100011010100100110000000001001000101010001110100100010101100111101010100110011100010000000000001000000000011111000;
    assign test_vec[39] = 1024'b1101100100011001010101011010001000010101110010110001010110000110000100101001011100110001000111100010010000100011100000100001110000000000000001100000100000001110001000001011010111100010000010110000011000001111101010101000001011111010101101110101001011000100001110001100001100001000010110011100011001010001101011000001000100000011110001100001010110011000010100010111000100000000110100101010011000100010101010011000010001110001111110101010001001010100001100101000001011000111000001000001100110110001010100011000111001000111111010110101000001010011000001001000100011100100010000001001010100101100111100011100011101000000010000110100100100000100000000010010100100111001010100100010000100011110001010100000010010101000001000010111001001001000010101011101011000010111010110100010100100001101101010100001000000111101000100100000001001111001011001111000000110000111001000000011000010010000010011000011010011100101101100001010010010010000000011010011000000001001001000000111011101110010101111000110000101110000001010000011001100110110;
    assign test_vec[40] = 1024'b0010010001000001110000011100000100000010000000100100101101010011010111101001100010001100001110100001011011100101000110001000001001101110111010000001101011010000011000000010001000000111000001111001010100100000000010001001100110111111001111010011000101010100011011001101001100100111101101000101100000011001001011011110000000000001100010100101000100000000010110001110001010001101001101010000011000100010100010001000000110000010011000110100001000000100010011100100111010100100100111000010100011100111000000000000010010010010110111100000000111010000111111010111111101010010110110101011010100000011100111010100001010000000111110011000101000011000111000101011000110010110111001101000100110001100000000110110110010101100001101011000100010010001100100111000110101110000010010001110010000011000100010000001001110100100001001101001111010010000000100100000001100000101010001001010111111111110110000101000001000000101000111000111111001111010000111101000100011000011010100000001011000000000101001100000011000101010100001000001100111100110;
    assign test_vec[41] = 1024'b0001000111110000010111100010111100001000100101100011010000111001011111100000100101010100111001000001111100010100010100000000000111011010101011000010000101110001000000011111101000100000010001001110010111011010011000000100010101001100111010000101100111001001100001001000100110000000110111001000001010000100010000000000011010100001000100100111110110001011001101011000001000000100001101100000001010111010010000001000100011100011011000000010000010110001011100010011000101000010011000010100000101101001001010011100101010001001110010111110001100000110000011010011111001000000111110010001100101100101010011000111010000000101010001110100101000111010010100010100100010101001110101001010110001101000110010010100100100001011010100000010101001001111011000011110001000010010010110011000011101100000001110000101001111000011110001100010000011010000110110001110000101011100110111101101010000111100000110110010101111010010000000001011010000110011110100111101000001001010011100001010100100010010100001000110001100100001001100000001011111101101;
    assign test_vec[42] = 1024'b0111000110001000011001010011101000010010000001000110001001100000000110111011011011101011100000000010010111111010010000010000101001000000101101010010110111110100011010011111110001000100010000001001010100111100001001011000011001000011001010011110101100010101100100111011000101110100101111010110110000000100101000100100010011101101010010000010000011100010110100001001101010110011001001000101100101001011001010000001011010000011001111010100010100011100000001000011010101000000011010010011010000100100000010100111110001100000100011000010100100101111000111101110001010011000001101000010011110000000010010001000100010111000011011101000101000010010111001001010000011010001001101011011100100001000110001011001101010001101110101011000000101110010110010011101000101101101000010010100010111110000111000001000001110010001100000000000100111010001100001110010000101010010110011110001001000000011001101010001101011101000010100100001010010001001110011110001110101000000101111000011011011101001001110101101110011110000000100011111111100010000;
    assign test_vec[43] = 1024'b0010111100011010010010000000000010011110000111001100010000100110001000110111011011100010010101000000000011010001010111101110000111111010110000000010000001010010101100011100110001110010010110010101100110110001100001010000100100111101111100000100101110010011000001000000010010011000010100000101110111111100010000111010100010100111110100010101101110100010101010010100110011111011011000100101001000000001000010100101011000011110100110001000000000111111100001110101010001011011110000000111011001000011011100101110001111000001110000100000110101010110100100101011010110000000010101000000110000100100001101000000010101011101000001011011011110000110100101101100010100000011011110110001010111111010101100100000001001100000010011000111001110100110011111011101101101100101001010100011111101100111110011010010010101000000000101000001100000000010011101011110110001100101100100001101101110100010110000100000101100100101000111110100101000011101000000100100010100001110101011000011100100011010000111100000100110110000010001100010000001000010;
    assign test_vec[44] = 1024'b1101100011011000100001110110111010000001001011010000100000111110101001011111011001100001010110110111010101011101110011001001001110101101011001011001010001000110000001100000111100110110111000000100001111000100100110001000001000010110000101100101001000000100100010000000110000010000011110011001000111001100110100100010101110101101101011001100001101101001100110001101101111011100110101110010110010101100111010100000111000001110110010000101011010111010011000000000101010100111100010110000001000101100011000110111001010110111011101110100001010001100010111010001010110000111101101100001101110001111000100000001011000010000000100000011110011000010100001101011010000100010101000011001100001100011000000000001000010100100100000101000101101000001000001000100010001110110011111011010000001101111011011110001100101101000001110101110010110100101111001001101001000000101010111111110110101000111100100101001001001001000011010001001010101001110110001010001001000000001010100001111100100110100000001001001011000100100111101010110010111010011;
    assign test_vec[45] = 1024'b1100111100110110000111101000000111100010001010000111101101000010100001111001100111010011011101110000101001010001001000001101110001010000101100101011110110001001001001010010100110100111001110101101000010001101100110001010110011000110011011111010110000110100110101001100001011111010101001010001100000110110101100010000010110100011101100111110110000111001001001000100100110001010010011001101011000101100010101000001001111011101010010101100010011101111101110001110001101001101001000011000010001010001101111110001001001111111110001110001000000110100011100011010010000101010100110011100011001101001111010001000001001110010100101110110110001001101001001000001001110100011001011010111000110010000000100101011101101000001111100000010111010100001110110010001011000001100111110001000000000010010000001100110101001000111001100001101101000000100101010111110100110100001110011001010100111000100010110101010110000010000101010111010100100001001000110100101101000001010010010001001010001110011010000010000000101001000011100001101110001111110;
    assign test_vec[46] = 1024'b1100110111001010101010010001000101100011000000010000110000011010010011000110011100010101111010000001000000010111011100010000011100111100000001010000101000000110000110010001110110000100111100000100000100000111001101001001110101110000111000100011101001011101100000000001010010100101010100010101110000111110001100001100011000110001001110000101100111100100110000000101001100101111111010111101111010100100000101001011010100011011010011001010101001100010100011011010110110110011010000000010111110101010001100010110001100101001100110100100011110110001011011100001110001110111001001100011111101010011100010000111011010000011100001010110010000010010101001101111001111111000000001001000101101000000000100111001010001011111010101111001101110110101001011100110100010000110010100111010100000011100000110001010101001001101111001101000111000010011100111011110100100111000111011100101100100111110001011001111110100000011111110010111001011001000001101111101111010000100111110100110000111000110000100000110110100001011011011100100011010010011;
    assign test_vec[47] = 1024'b1011110011101000011011011101001110111101010001010101100000000100100111000001100010110010101110101000000111001000101100001100001110000101011001110110110001000010011101100000111011100100110001001001100011010001000100111001010111110000000001101100010000110111100001110000000010101100011101010000101110011110110001010101001110110010010011011111100100011000010011011110000110001010110011000011100100010010000100010010011010111000101001011100100000111111011100101000100000111000100101110100000101011100111011101001000111101101000001000111110001100100100110001110010110001110111000001001111100111110001010100000100000101101101000010100101001011000100110000000101100110010100000100000011110110001101101011011100111111011000000010110101111001010001011001101111111001001000100011100010010010100001101010111111001101001101000101110001011011100011101011101001101110001001011010010000000010110110111110110100010101110001011000111000111010100100000010001110101001000011001111001101011001111100111101000011011100001100011111011110000101101;
    assign test_vec[48] = 1024'b0010001010100000001110001001100011110011010001011011111101100111001000101111001010010111010111001010101000000010010101001010000110100011011101110001001111001111010101001010100000110000111000111001100100000110110010010010001110001101010110000110011000110001110010001011010101011001010000101000111000010010111110001011111011001110110001101111101010101000110110001001010010111101011101101001001000000100001000011100101010100011000100110011110110111100111011100100000011001010111001001011010010110101010001011101011011100101111111000101011011111111101010110110001010100101111111010100000001100000000110100010000010100011011010111001100110001010010011110111001110100110011100111110000000100111101101100010111001101001110011111000001100010011001011110001011110110000000000000001110101010100011000010011000101100000011011000001101000000000000111101001100010100100010101011111011110001000011101111110100110101000100100011000101111110100001011111101011001101101110000001001111111010100011000101011001000101101001000100110011101110001;
    assign test_vec[49] = 1024'b1000011010110111110001110001111101111010111101010110101000110111000100001101101000110110111010101000101001011110000101011001001001110010100011010001010010101011001110010110100001100001001001100000101011011010100011010001000110110000000010111100010100101010101100110101010000110011010011001010110101000110011100101110000111001110111001000011111011110111110111011010010000100111110000001000010101011010011001001100010010011011101010111001101011100110110010100101001111001110100111010100000100001111001000101111100000100101011111000011010010000000101100101110100111100101000100011111100000010111100101000111001101010010001000100100001111001110001010000001010111010001010100010111010100101001010111101100010101110101011111100110000011001111110110000101011101101110111001101100100010101111111011010010011100000110101001010100100110101000011100101011001100101011000011001110000111101000001100001101111011000001111111010010110010100111011001110110101100111011100110000000110001101000000000110010001110001100101010101011000011111010;
    assign test_vec[50] = 1024'b1110001011000111111001000100101111101010110111101011000111100101111011011001111100010011000101011111110010000111110011011110100011101111101010010010000001111110001110111111011100111101101000001100100011001111100100010001100010111011010100001001111111101001100101010100001011101010111100110110000001101110111000011010000101001011110111010111000000000100111111111001100100000000000100000100100100100101011111001011010001101001011000000100100110000111001011111110001100101000000000101010110000111010101010100110010110111101001110000101010110011010011000000101011010111000000001100001110100101011111010011101110010100001000100010001001010100001110110101100100011101100001010100010101111010011100010011100111000110011011001100001111011111101000011010010101001001111001110011100011011011101110110110111011100101010100010001111100101100011001110001001010011111011111110001100100001011010001110000011000011110111101110101101100000000111101110100100110000011110111100011001000110111000100001010000100010010000011001001110010110110011;
    assign test_vec[51] = 1024'b1000000111110011010101001011111100000010110001011101010101101000010001110001011110101000101100000111111111010111001000010011001011011111111111011001101111111101100110001100100100111010110101101111001100011001111101000000001011000000001110000000110011100010110011000001101111011100000000000010101010011001000110011001100101010011011010011100100110010100111010100101000000000100000100010110110011101011111101011001110001000001011010101111101100111111100000001010100101011100110101001000110011111001001011111101111010001111101001000010101011110111101100111000010001010110110101111111110011101101001110111101101000001010000000010000010001100000001100111010010000010111111010110000100011101110101101011111100111000000100100001101010010111101001111110111110001010111111101001110010010010101111000111000111110000111101010010111011101110101011010100001010110110001010110110001011110100110100001001101011111100001100101101011101010101111001100001001011001110110111001100000010100000000010111100101000100011011111110111010111000011011;
    assign test_vec[52] = 1024'b1001111100100111001001100010101000010111001111100001101011101100010001111011110111110010001111111010100011010110100111011111011110000011111110111101110000110001000100100001111101001100011101111110111010100001111111001101001001010101000011111111100001100010010111010001000011110101100001011100101111100110110100011110101101001011001111011011000100000100000010000011011110110100000111110110000011011100110001111010101111111110111111100111101000000001111110100110000100111011100011110110100101001011000010000111010100010000000010111101110011100100010001001000000111001100111001101011110100110011111111100000110000111001000000001100101010011100011110001110101001100010001111110111000101110111010010001111101011010001110010011001010000111010100011101001100011100101011111001110000010100011110101000111101010000101100101001001000000000111100111101100111001011100101010011010111101111111100000000011001010001011010000110011111000100001011010001001000010011011101011101110010000110111010111011111001101111110000110001111111001101001;
    assign test_vec[53] = 1024'b1100111111100010011101111001010010000011111000010110011110000011010001100110110001100011011000111000101110111001000000101101111110111001000100001111110011100100110110011010001011100111110001001110101110000011111111111001011011011111001001101110111101010010011101101101001001010011010110011001000101100001101111011111000111111110100111011101011001010010100111111011101001110011100001010110010000101000110100011101000101000111010100110001111100000100010101011011100111100101001000001000101010111110110001101110010001101000110111011011110111011101001001001000011011100101110111000111001111001001001001101000010111110011101110001001111101101110010000000010001110011000111000010111010100011101101010100100011000001000000111110110001101001101111111011000110011101000001111110011001001111100010011110101011001111111000111000000011010110100001100100100111101101111010100110101111100111110101110001100001110111010011001100010111101010100011110110100101011000111011110000111010100000110101110110000100101110100011100111101001000110011;
    assign test_vec[54] = 1024'b0010100011101001011001111111100111101001101110010010111000110101111011110111000000111111100001001111111011100001111001111001111011101001101110110001101010011111111011011111110101111010111110110110110010111111010110110111110011000100100111000010011100000011011010101111010000100111100001001110100001001001110000110011110111000101001011001100101001111110110010000101100010010000111010000010010111111001010101011001101101011011110101100100010111101000011110010001010010111101100011101110101100010111010101111001111111101110110011111100110011001001001011010100111100010001110010111100101110001101111101111001100011101010011101001000001111101001110111000100110100101110001110100110111001111000100110011101110001000001101100011101110101001111101110011011110010000101010110001011001100001110111000100100100100001101101010111001100100100001001000001110100011110000000001010011000111001010000110011110100001111110010001101111010001101111100000010000001011001000101110110111101001111111011100110100001111111010001010001011100001110111;
    assign test_vec[55] = 1024'b0111011110110000010001010100111000011110011101001110111001000101011011100001110001001110111110100101001011110001100111101111111111111100011010111111001001011100111100111110111111000011110111000100010100000111011100011011000001001111101000101010000100001001110011001100100010001000101010000000011101101001001111111110110010011110011100100010111010010100101000011111000010001110011110001110111110011111101101011001111111101000101010000101011101111100010111011100110001101001101111110010011001101011011100100011110111110101011100111101111100111100101010101001010100101010101011000111000101001000011000111001111011010111011101010100100101011100110000110101111010101111111110111110010010011111001010101100010101100010010100111101011100001001010111000100100011111010111100100101001110001011010110111111110011101011000101001010101100010101001100110010101001111000010010110110010101110111111011111100011100111010011011111010100001100110111011001110000101000111001111110110110011001010100101111110111110110010000010100100111100110011;
    assign test_vec[56] = 1024'b1011100011111011011101101011100111101100000000110100010000100110000111111000110000011100010001010010010110100101101011001110100100111101110011101100011111101011011001101101101011010111101110100111101010101010111000010101111111101011001110010000100101101111001100011101100111010101011010101100100011010111011100111010111101001110001010101011011111001011111011110101100011110100100110010001000101011110111011011110101111011110100110111111111111000001101000111100011001110100001101000010101010011110001110101010110100111111000111101110111000011000010101000101100010111111011110001111100100000101010011111011111011101010101001111110011111010001111011110110110111101110000111000000000000000110100100101010111110011110111101101011101111011001010110100011011010011010001000101110000011010010101101111110100011010111100000011100010001010001111110000010110110110000100101110011101110011000001001000010011010110101110111000101111010110011110010110110101111011110110101010110011001011000111101111001100110101101101011001111111111011110;
    assign test_vec[57] = 1024'b0100100111011110011011011101101101110101010110111110101111011011101110011000011001010101110101001011100100100110101100001110001111111011100111101001001110100011000110011011011110111001100110101101000110000100110001111011011010110001001111110111101011001111101011111000110101011101001111110101111110111101101111101011010101001011010011000111101100011010101110111100100010101100110101010111101100100110100010001111101011111010000001001000010111110011100001110011000101110110111001000110010000110101010001010001000111101010010010110101111110111111111111101100111101101011101111111111011000011100111000011001100011110111110001111011100111011000111111011100100111110110011101101111011111011101001100001111010111001010011111111001001111000000100111001110110011100101100100101111101000000000010110011110111111010111111111100000001010111011000000000101110100111010110001011100110111100111000010011110110001010111010100111111011001011101110101011111001101000000110100101010000000111001111010011000101001111000011011000101100110011010;
    assign test_vec[58] = 1024'b1001100111111100110011110111011011001110101110111010010001000010010000011111101101010000001011001011101001111001111010111101000101000100101110101100111011110101010110001101110111011010011000111110001110001001011101010101111010110111101001101111010110110111111000001101110100110010010001011001110100011010101001010111111111110111110010111011110001111110110011101111011110111000001111011000011110000110110001111101111100011011110110101001110011110111100011101100001011110111101011111000001010100110000010111101101001111100110100101101110101010100100000100111100111101100100100010011111101001010000101111110111110010100101011101111000001011100011110011001101110010111011000001111100100001111000011110101001110100111101100010011110100001111110001101010010111010011011111001001010111010001101100110001001100101111101011100111111010111111110011101101100011111110111010011101010001011111101000110100101111010111110101001111111110100000001000010101111011101100000110000111110110100101110001111110010011101101110011101110111111100111;
    assign test_vec[59] = 1024'b0011100001110110001011010011011101000111010111111011111110110100000001110011011000001001110000110100110111111001011101111011111010011111000101001010000010001111010111101101100111110100111011011101001111011110010111110011110111011011110001001001110101010111011101110011011100111010101011111101001011000101101110011000101111010110101111110100011110101101111010100101000011101100011100010111111001111011001111100010010111010110011100111110111010110010110111111101001010110111010101101111001101101111010001010000100011010100100000111001111101111110110000011111110010101100011001010100100101110101011001001111101010111111110111101010101111001000001010110111010101100100111010001110101100010101100111111011010100001000111111110001110111000110010011011101110100011001110101011011111000011111111101110010110100100100101111111100011011101000001101111111111111000111011101000011100011111111110101110101001011101111100110000011111111011010111111111000111101001111100001010010110010110111111000110010011001001001111110101010000011010111;
    assign test_vec[60] = 1024'b0010111011111111000111100100110111101100110111110101000010011101110011001110011000100000010111101010011111111111100001110111110000010001101011111010011101010111101011101101001101110111111110101010111101111111101010010011110101001111110001011011111000011111011110000101001001010101101110101111110000100100010110000010101111111010111010100010110101001111000010110100011110111110001011010101111001011110111111101110101000010011110110001011111011010010110011110111111000011111011111111110011000000101111001101010001001110111110101101011111111100000100011000111111011101111110101010110110110101001001110111111100001111110011011101011000110010111110111111011100110011101111111101110010011001100001101101101011110111000011001101110111101111111000110110111110100010110111001101111000110100110111010101110000010110111101110111100100111000011110100101100100111011111001101110000010111111011111111001101100011001010101111011101010111001100111010100110100100100011111110000010011111001111010011100010000111011011010110101000101011101011;
    assign test_vec[61] = 1024'b1101111100100010110111001110011111100111111111011011101010111101111001111101111111111001101110111100111101110010101100110001101111111000001011000111101100010010010000011110100110111011111010010010010011001111101010011011001000101100001110100111011011111101010101011101100111101101111101000111011111011101101101111110010100010101001111010111001111111110010111111011101001111001010111110111010111001010111111011010110100100011010111111110111110011010001011111110111111100110010000110010100100111111011011011001110111100011011011110011111011010011111110110101001100000110001110100011011111011110110111011110000001001110110010010111001101111111111101001111010111101110011100110000101111101010111010110000111000011010100100111011100111110001110010001101101101110011111111101110001110111110110010100101110000011101110010110110101110011111100000101111111110101000011110110111110001011000110011011101111100001100101111110011101011001011100110011010011110111101010100110011111111001110011111110001010111011000001001010010110000100000;
    assign test_vec[62] = 1024'b1111110100111101011110110110100011011100001110011010111110111110101010111111011111110010101110110111001101011011110100111111111101000100100101011111100011111001110101111111111111001001110100100111111101110110101100110110001010011000110001010100001111111011100111001111111001110011101011110010111110001011110111011100101000111100110101010101111111111100111101011000011111011110100111010100111001101111100111101010111010110100010100111111011101100110110000011111111001000000111010000010111011111111110100100111000001000111011001100111110101101011000001110111101111100111100100001101111101000011111111010100010011001100000001111101011110111000000111101011000111010111101100111111111110001110011111111001111101001100111101110011100101110010111101110011100100101001000110010111101111001010111011100100111110110000111001011101001010010001011111101001111011011011111100111010111111101010000111011011001111110100111101001111010010111011101110101010111111110000111010101101011110101011111101111101001100101011110011010111101110101101;
    assign test_vec[63] = 1024'b0100000011111100010111101101101010011001111000011101100101010100110111010011001011111110010110111011101011001001111111111011111100111010111101001011001001111101110101111111111111101101011010000110011101111001101101111101001110000111110000111110001111100011111100101011000101111001111110011111101000100101110011111101010111101111111111100111101001111111011010110101010001110111101101111111001001011110111101001101111100101001111001111101101111010101011111110110111111111111110111101011011010111101011101001111110111001101111001000111111011011111100101010111110111111111111100010011111110101000011111010110110101101000010111000101000010101111101011111111001101101011001100111101100111100001111111111011100111000000111011010100100101111100010100011111111010011011001010000100011000111001111001111100111100001101101101011101000111111111101101111100011100000100100011110110111011010111011100011011011111110111101001110111110000101000101001111111001101010100011010110011010101111010100111001010011101000111010101111111110101111000;
    assign test_vec[64] = 1024'b1001111010101111011011110110010101111011101111111100101001101101001111101111110110111100111000011001011110101110111111011011010000111111001100011101101111010111110001001111011110111111110110000111101111011111110011110101001110011110011101100100011110111011111011011001011011101111101110111010111111110010111111011100111101010111110100110010001111111001110101110111111110101010111110101111011010110010100101101001111111110010111001110110010110110010001010011001101010111011110111101110101111010101110000010011101011110111010001010001111000101011111001100110011001111110011111110111100001101110011010100001111000110011000111010111101001110001011111111100110101110111111011001110010001110010001011101111011100101011110011011010111111101011011101001111111111000101011011001101110110111010110111111110101100101110111100011111010011100010101111110110100111011111111011111110011010000110110011010011101111000010010110111010011110010110110000111110011011111010101111100011110111001011010100001110111100011010011101110101011111110111;
    assign test_vec[65] = 1024'b0110101111011010110001010010110010111111110111101011010111000110000011111011111100100010111000111111101001001010010111101111111011110101110110011100110111110010101111100111101011110101011001110111011101100111111111111001111111010001111001111111000101111101011011001111001110111111110110000111101111111011011011111011111111111101101101111111100100001000111010111110111011001110101111010110101101101011111101101010000010011110110111011000110101111100110100111011111000111111111111111111111001111110111111010111110101001111001110111111001010011011111100101101101011010000100111110001111101011110111111110111000011011001100100011110011000111111000111111111110011011010110010111010101101001010101000011100001100111010110101110010001100111100010101001101111101011100001101111101110111011100011111111110111111101011011011001110011011100110011001101111100001010101111110101011001101100111101111001011001110101011110001101111110011110111111010011001010111001011010100110000101010111111111100110110111111011101100001111111011011110111;
    assign test_vec[66] = 1024'b1010111001111111111111111110011100011011100011111110001001011100111100110010110101111100101101110111101110111100100011111011111101001110111100110001011110111111101001011101111110011001111111010101101101111111011010101100011110000011010011011001011111011011010101111100111100111101000011111111100101000111111000011111101100010111111001110110111011100001111110110111011111000111110011111100111110100111011111111010111101111111110001010111111010101111110011100011100110111101110011111100111100001101111111111100001001001101111011101001110111010100110111111111110101011011011101001101001101111110111111101111110100010110110110000101000110110111111101100001000111011000011011001001101001111110111001111101011110111101110110011111111110111001001100110111001110110011111001011011000010011110111111111100110000011101011000001110001111101000011110011111101111110001010011010001110101011000100110101010100111101111111111111111101101111110011010011001111111111111011111111011100110111110011001010111111111001101111001110111111001111111;
    assign test_vec[67] = 1024'b0011010011001011110001010010011111101011110100000110111110010101011111110101001011101101011110110100011111111001110110011011110111101111110001111110100111101001101111010110100100111111101001111011101011111011110011111100111001101110101000110101111111111100101111111101110011110000001111011111110100000101111101111101111111010111011111100101111100101110110111011101111111101011101100101111101001010111111111011111101111101010111111111011100011000011111111111001001101011011011101111111111111001101101000011001011101110101101101111010110100111011100001101101111001010111110101011101011110001111111101011111111111101010111101110111011011011011100011001111111000101101000111111110100111111111110110011000101111011101111011101010011111010011101001111110110001111111100101111000011111001010110011000111010000110110100011110111011011011011011011011001001010101111110101111110111111101111010101101110111001101101111111110111010011111010111111111101011010101101011001001100110111111111011001111110111000111110101100011111011101100111;
    assign test_vec[68] = 1024'b1111100011011100111111111110010111111111111101100011001111110111011111111100110111001000011111111011000110111011101101011011111101010100000101100111101111001111011010101111101111001001110011010111101101001011110111011111011010011101111111101111111111111101111100111011111001100010010010111001011000110111010111011100100000011011111000111111110001111110001101110011100001101111110011110111101101110011111110111111111101101110101110101101011111011001011111100100101111111101011001101011111011111101101101001011100101111110111111011111011111111111111011100011010010111101010000111000110111011111011011111011110111111111111101110111001001111110011011111110110110110111100100100001011100110110111101001110111101110001111111111111011101000111101111111011100110000010111000111000111101010110111111110010110111110101101111110111110111011111110101011000000111111100111111111011011111111110101110111110101101001100011111100110111100111011111000100011110111011111100101101111010011001101111001101110101001110011100100011110011101101111;
    assign test_vec[69] = 1024'b1010111011101111111111111000000111001111111101111001001110011111101111110101011111110010011001110011100110000100101011011111011111000111011101011000011111001111111111101110111111010011111101111011111010011110000011110101111101011110101011100001110101111000011111110011011011011011011101111111111000000111101111010011111111100111001101010001000101101101110110111101101001111111111111111101101110110011101110111101111111000011101011101011101100110101111100111111110001111100111111011011111111111111101000100011110111101110111100101110101000110100111111100111010011111101110001111110111100111110011111010011100101111011111010100101110110111010001111110100101011111111101101110001011011101111111010001111111111010111101001111111111111110111110011111101010010110111111111001011111111111101011100010111110001111101000001011111111011001001110101110110011111111111110101111011010110111101110101101100110111111100110000100111001111111011111011111111101011101111000111011101010110111011110011010111011111111111101110011111111111010010;
    assign test_vec[70] = 1024'b1010011100011111011001011111111110111010100011010001101100100100111111110111110101111001011110111111111111111101011111000110101010101110010011111111101011101011001001011111011011001111101111111100010111111100101111100110111100111110111110110110101011110110111001100111101011011111110110011111111110110000010101111111110111110110101101101110010100111111111110100101011001001111111001101111110111111000010001111011010111011000111111111111011000110010011100111101111110111101010010010111111010011100100100111101110111011111111111011111111011010101110111100111011111001101111011111000011011110101111111111011110110101111011110111110101101010111100111110101011111111111011001111101111100111110100011010111111111110011110110111110110110110111111101001111111111101010111111100111111011101101010111010110110111111010110011011011101110011111000110110111001111001011011011111011110111110111001011101111111110111101101111101000010110101110110111110101111100111110011101110101111111111111101111000101101011111111011011110111011001011001;
    assign test_vec[71] = 1024'b0111011111101100101100001111111110111101101110001001110011111110011011101111101010111010101100111111100111100101001100110101011101100011001011111111100101111101111111100001011101101110111000110101111111111000101011101110111110010001110111010111110100111111111111010101111101001110011111110101111011011110110111101011111111101111111110011110111111110111011100111001111111101011110011111100111001101111110111100011100111111011111011110011111011000110111011111011111011111011001111011110011011111111011111100000110111111000111011010011111001111111110101011110100110111101100110011010111111101010110111111001101111110100010010110101110111111101111111011011001111010111111111010111100111100101010111111111111111011111011011101110101111110101111100110101111110110111111001111011111001111111011111110010101011010010111010110111111001110101111011011101011111111110010100100111101111001110111111101101110111110011011111101111101111101111101001010111111101111000111111111001010111101101110101111110011110010111101110111111011001111011;
    assign test_vec[72] = 1024'b0101100010101111101101010001011010111111001101010101000111111111111111101101011110100100011010101010111111111011101001010111111101101000111111101011111011010110101000110010111101111011011111111011110100101101011101101011011111111111101111101111111110111111011111111101011101111000110100100010111001111101011010111111100111111111100110011111110111010111101111011100101011111111111110101101110111011111101110101011110000111111110011100110110111101010111100101111011110110101110000111001011111111111101111111101101110110101100111011101111101111111011101111111001101110110000011111011111101100111010001101011010111111111011011001110110111101100111111101111111111110111111101111011100111010111111001110111101111111111011000110111111111001011111110110111110011110111111111110011000111011101110110111011111011111111111010110010110001101111110111001111011001111001110011101111001111110101101111100011101111111000101101011111111011110011101111001111010011111111111100101011001111111111111111101111111111011101101111111111111111001101;
    assign test_vec[73] = 1024'b1010011111000111101101011110111010001110011111111001110001100111101101110111111011111111110111111111110111010101110001111111111111000111110111101010110110110110011110011001101010111101111011011110110010101101110111101000011111111101100111001111101111111111111010111011011101111110111111111011111110101111111011111101101010101011101111011111110110111001111001111111101110111011110101110010110101100110111111111001111011111111111011101101110110100101100110101110111111110101101011111111010101011111101111110110111010101010010101111010011001011100111100111111010111111111111011110111110110001011111000111011111111011100111111110111100111010101110011001111111101110111001111100111111100111101101100111011011011111111111111110111110101111101011101111111110011111110001111111001011011111011101101111110011101001101101111111101111101111111111101111011100101001101111101101111011100111011001011101111110110110101111001111111111111111011101000011111111111111101011111111111110110001111111011110101111011101011111101011110001010101100;
    assign test_vec[74] = 1024'b0110001111111111111110111111011111011011101010001111111100110110111111101111110100101011110111101111110111111001100111111011011111111111001001101011000110011110111001111011111011110110111100111111101111011011100111010111001011101101111111011111111111101110110101011111001000110111110111011111111111111111101111010110110111111111110111101001110110111011111111100111111111111101010010110111101111111111111110101111011010011111101101110111101100011111100011010110011110010111111001010111000110101001111011011000100110111110110111111111111111111111111111110111011111101111111101011111111011111111111010111111011110111011111001101101010110111111101111111011011011000101101111101101111111110010111001011111011110110111010111011101100111111011011111111011000100000111101111011100011111111010101111111111110111011011111000001110001001101100111111111111110111111111111110011011110110111111110011011101111101111110111101101110011111011111101101101011111100001100111000111111110111110110110111011111010111111111010101101010110110111111;
    assign test_vec[75] = 1024'b1101111011011111011111110111111011111111011111111001110001101011110101111111011111111111111011101110100011010001111111111110011011100011011110111010100100111111101111111111111110100110111110100111001111111111111111111111101101111011001110110000010011110111011111111111111101101111101000100011001101011110011111110100101101110001110101010001011111101010111111110011111011111110011111011110011011110101100100111111111001111110111110110111001111011101011011111111111101011110110110011111111110111101111011101001011110010111111101110011111111111111111111111101111111100111010101111100101011101111100111111111100011001111000011011011111011111111111111101111111001111111101101011111110111110111101100011010011111101111111011101110110101111001111111111011110011111111101111111110011111111100111111111011111111110111101111101011110111101111110111111111111010111101011101111101011011110111010111101111111011011111101101111111100111111111111100110111001011001011101111111100101111111111111100000010111010011101101011110110111101110111;
    assign test_vec[76] = 1024'b0111001111111011111100010111001111011111010011111111111111111111111111011010111111001111011010100110011111101110001110100111111111100111001011100110101101100010011011101111110111001110000111011000011101110101111011110100111010110011111111111110100001100111011111111101111011001010011101111111111111101110111100101111101110111111011111110111010010111110111101111111101111011101010101111111111111011011111101001111111110111011111111011010101011101011100010011111111110011101110111111111111110101111001111010011111011111111111111011110100011110100110010111111111111111111111110111111111111111101100111110011111011011111111111101111111101111110111110111111111111011111001011110101111111111101111110011101101111111111110111100011011111111111101110000101111101010111001101111111011111001101011110111111111111111111011110111011101111111111111111111111101111111001011101110101100110110111101111110111110111111011111111101010111011111011111101101001101011110101011101110110111010111100101011101111111101101111010111111101111111111111;
    assign test_vec[77] = 1024'b1111111111110111111011111011111011010111111111111101011100011111110101111011101011101111111111001110011111111101001111111110111110011001111101100101111101101110101010111011001111011110111110000101111111011101011110001111111001111111111111011111110101111111110111111111011111111110111101101110111111100111110111011111011011110111010111111111101011111000011110101111110110111111111111101111111110111111111011101001111111111111111011001110111011011101101010110111110111111110110011111100111111101111110000111110111111110111111001101111111111111111111101111111111011011111011111100111111110111111111111111101110010110110011111100111111111101011111101110011111100011111010111001011111111011011111111100101111001011010010110101101111111011001101111111011111001101110011110111001111110110110111000110111111100110101111010110101111011111111101111111011101010111111111111101111001111110011111001010111111101001111010111111110111111001111110101101100101111100100111111111110111111111011111111111111100010100011111111011111101101111110;
    assign test_vec[78] = 1024'b0111111101111111011001111101110001111110010110111101110111101111110101111111111001101011011010011110111111110011111010111111011111111111011111111001011101110111010111111110101111101111111111010100110101111000111111101001111110111010011111001110011101111011111111111001111010011111110111011101111111111111110110101111101111111101111111010111111011100111111110111011111000011111011110011101111111111110111111111111111111101111111011111111001011111111111111111011111100110111011111101110110111111101111111111011111111110110111111111111001111101101111111111111111011011100110011011101010111111101011111011111100110110111011011111111011111010111001111101001011101110111111111010111110111111011011011110111111110010001110111011110101011111111011011001111111111110111101111110101111111110111111101111011110111111011111011111101010011111101111111100100011111100011010101101111111111101110100001111011111101111001111111111111111000111011011111111111111111000110111111111010011111011110110111110110111111100111110101001111111111111111;
    assign test_vec[79] = 1024'b1110111111011111101110111111111111111111111111101111110110111111111111110010101111011011101111110110100011101011111111111110111111110101110111111110011101111011111111101011111110111110001111101001110111101101110111110111111110011110110011111111101111101111000110111111111111011111110100111111111111011010101111111111111111101101011011111011111111011110111111111101100111011101010111111001111110001101110111111111111010111010111011111111111111111111000101111110111011101111110111011011011111011101111111111001111011101111101101101111110110010101101111101111111110000011010001111001111111111111101011111110111111111110111110111001111111101111101111111110101111110110110001110111011111011111111011011101111111011111111101101101110110111111111101111111111100110111110111011111111111111011110111011111101111100111000111010101011110111101011111111011111111111110101111111011111110011111011111101111111111011111100111011111111011111110010010110101011111010011101111100101111011011111000111111111111111001011110110111101111111110111;
    assign test_vec[80] = 1024'b1111111010111110011111111111011101110111111001011001110111101111111111111010011110111111111101111111011000111111011111111101111111111110111011111111111101100111110111001010111111111101111010111111111111010111111001111111111001011111111111011011111110111011111111111111111001111110111110110101011101110111101011001011101011111110101111011101101011111100110111111111101110111010111011110111111111101111111001110111111111111011111111111011111101110110011011011110111111111110101111101101111101011011111011111111111100111011111111011101111111111111111111111111110111001011111101111101100111011100111111111101110011111011111110110011101110111110111111111111011111100111111110111111001110001111111010110111111011111101101111111111111111011111111111001111011110101011001111011111011101001111101111111111111111111011100100110111101110111101111111010011111111111110110111111111101101111111011000111101111111011011111110111111111101100111110101111111011111111101101110111110111111111111110011111111000101111111011101011001111101001111;
    assign test_vec[81] = 1024'b1111001011100011111111110111011010111001111111110111111111101100111101111101011111101111111101111101101101101111111111111101101101101111110111111110011110101100111011111111111111111111110000111011111101111111110111111111110111100111111101111101110011101101101111111101100011110111111111011011111111110011111111011100111101111110111011010011111011111110111111111111111011011111111111111110111011111010111111111101111111111101111101111111111110110111011111111111110111011111110101110110111111110111111111110011010111110101011111111011111110110100101111110110111001000111100111111110111110110110111111111111111111111111011111011111011111111111111111101110111111101111111100110111011111111111111111111111111011111101001101111111111110101011010101111111111110111111101111111111111101011111010111010111011101110110110100010110011111111011110111111101011111111111101111111111111111011110111101101110011011011101111101111111101010011111111111111111111111011111111011111011111111111101011111111011110010111001111111001111011010101111;
    assign test_vec[82] = 1024'b1011111111011110111011111111111111011111101110111011111110011111111111111111111101101111111010110111110111011010111111100111111111010110110111000110111010011111011111111110110111111111111111111110111101101011011101011011111111111111011101010011111111101101111101111001111111111110110111111111111101111110111111110101110110111111111111111111111111010111110111111111101011111111111000111111001111110111110101011100110111111101111111011101101111101111001111111111101011110111101111111111110100111101111101110111011111110110111111110111111111111101001111111111101101111111000011111101110111111111011111100110111111110010001111111000111100001111110111110110111111111111111111111111111011111101110110100111101111101111011101011101111111011111111111111111111111111111110101011100111111111111111101111111111011110111011110111001101111011111111011111111111111011100101111101111011010100111111111111111111011111101011101101111111111110111011011011101011111111111111101111111111111111111100111101111111011111110111111011111111111111111;
    assign test_vec[83] = 1024'b0110101010110111111111111111111110111111111100001111111101111111111111111110111111101111011111011111111111001011111110101101111110101010111111011111101110101111111111111111111111111101111110111110110111111111111111111110111011011111111111111111101111010111111111111111111011111100111111111100110111111111110111101111111111111011111110000110111011111111000111111111111101100111111010111011110011110111011111111110111111111011101010111111101111111111111101111011111111110011101111011011011111111111001111111100111111111111111100111110111111111110110111111111111011111101111011111111111111001111111111101111111111111111111001101101111111110000111110000110111011101111111100111011111011111111111111111111011001110011111011111011011010011110111110111110011111111110111111101100101111011111011111110010111011111101111111111111011111100111011011111110110111111111111111001100011111111010111111011011111111111101111111111010111111101111111110111111110111111101111111111111011111111011111111111000011110111111011111111111111111101111;
    assign test_vec[84] = 1024'b1100111111111101101111110001101111110111111110111011111100111011111111111111111111111111111101111110101111111111010111111111101111010111000011111111111111111101111111111111111111111110111111101101111111111101101101001111111010111111111101101101011111111101111111111011110111110111011111111111110001111110111110111111101110111110111001111111110111111100000111011011011111111100111110111111101110111110111111111111111001111011111111100111101110111110111111010111111101111110111111110111110111111011111011101101111011111111011111111101011111111110111111111111110111111100101111010111110111111111101111110111111111111101110111111111111011111110111011010010110011111101011111101111111011011111111111111111111110110011111111111111111111111111111011000010100100111111111111011111111111011111111111111111111111001111111111111111111111111111111111011111110111111011001110111110111111001011111011111111111111111111001111011100111111111111111110111101111111110111111111111111111111111111111100111111101111011110111101111101011111111101;
    assign test_vec[85] = 1024'b1110111111110111010111111111110110111111111111010111111111111111011111101111111111111101111110111111101111111111111110111101011011111111011111111011111111111100100011001101110010110110111111101111111111011111111110110001111111111011111111111001111111111111111111111111111111111011011101011111110111111110100111111111111111111111110111111111111111111111111111111101111110110111111111110111010111110111101101111111111111010001111101111111101110110110110101101111101111111111101111111100111111101011110110010101111100111111111111110011111101110111111111111110101011111110111111111111111111111101111101111011111111111111111111111111101111110101101111111111111111111111111111101111111110001111111111111111111111111111111111100011011110100101111100111111111111110101101111111111110011111111111110011110101111111101011110111011110111111111111110011111111110011111111111111111111111111111111111111111110111111100110111111110111100111101101101111110111011110011111111011111111011001101111101111111101111111111111111011111111011111111;
    assign test_vec[86] = 1024'b1111001111111011111101111111111100111111111111111101110111111111100111011111111111101111010101111111111101101111111011111111111111101111111001101010101111111111111111111010111111111101110111111111111111111110111111111111111110111010111110111111111110111111111100111111111111111111100111111111011111111100101111110111011111011101011111011110111111111101111111111001010111111101011111100111111111110111111011111111111100111111011111111111111111111111011111111111111111011111011111111111111101011111111111101001011011111111011111101101111111111011111110011101101111111111111111111111111111101111111111111111100110111111111111111110111010100110101111111011111110011111110111111110111111111111111111111111010111110111011111101011010111011111111111011111111011111111111111101111101111111011111101110101111111111111111111111111111101111101111101111111110111001111110011111111101111101111110111110111111011111110111111111101111000001101111111111111111111111110111111111101111111101111111111111111110111111111101111111111111111100011;
    assign test_vec[87] = 1024'b1111101101111111111111101110111011010111110111111111110011011101111111110111110111111111111111111111010111111111111111111111111001111111111111111011111110111011101111111110110110111110110111111101111011011110101111111101111101111111111111111111111110110111101111111101111110111011111111111111111101111111011010111111111111111111111111101111111111111011111001111001111111111110000111111101111111110111010101111110111111111111111011111011101111010110110101111111111101111011010111011111111101011111111111101111111111011111111111111111111111111111111011111011111111111011111111111111111111111101111011111111111111111111110111110101101111111011111111101111111011011111111111111111101111101101111111011110110111011111111111111111111011111111001111111101111111111111111111111110111111111110110111111111101111111001111111111011111111111111100110110111110111111111011001101100111111111111111111111111111111111111011111011110111111111111110111111111011111111111111111110011111011111111111111111111100111111110111111011110110111111011;
    assign test_vec[88] = 1024'b0101111011011111111111011111111111110111111111110101101101111110110111111110110111111111111101111111101111111111110110111100111111111111111111111111111111110011111111111111111010111111111111011111111011111111101111111001111110011111111011111111111111110111111111111110110111101111111111111111111111111111111111111011111111111111111111111111111111001001011011111111111111111111110111011111111111111111111001111111111110111111111011111101111111111110110111111110011111111101101111111111110111111101111111111111011110111101010011111001111111111111110111111111111111111110111111111111111111111111101111111101011101111110111111011111111111111011111111111111111111111111101111111011111101011111111111110110111101111110111111111111111111110110011101111111111011100101111111111101111111111111111111111110111111111111111110111111111111111111111011111011111111111111111100111111111111111111111001110111111011111011110111111110101111101100110111111111111111101111111110111101011101111110110111111101101101111111111111111110111110111101;
    assign test_vec[89] = 1024'b1111011111111111011111111111111111111111011011111111110110111111111111001110111111110111110111111111111111111111111110111111111111111110111111111110111111111111111111111111111111110111101101111111111111111111101111011111111110110111101111111111101111111110111101111101111111110111110111010111111111110011111100111111111111111011111111111111111111111111101111111111111111111111111111101110111110111111111011111111011111111111111111111111111110110101101110111011111111011111111111111001111111111110111011111001111111111111010111111111111100111111010101111111111111111111111101101101111110111100111011111111111111111111111111110111101111011111111111011111101011101101011111111111111111111111111111111111011111100111101111111111111111111011101111111111111101111111111111111001111101101111111111111111111101110111101110111111101101111111101111011111011111111111111011111111111111111110110111111111101111111111111111011111111110110111111111111111011011111111111111111111111111111111111111111111111101111011111111010111110110101111;
    assign test_vec[90] = 1024'b1111111110111111111111110111111011111110011011011111111111111111111111101111011111101111111111111111111111111111111011111111111110111111111011011111111111111111110111110011111111111111111101111010111111111111101101111011111111111110111111111111111111111111111111111111101111111111111111111011111111111101111101111111101111111111111111011111011111111111111111111111100110101110111101111111111110111111011111111111101111111111111001111011111111101110011111111111111110111101111111101101111111111111111011111110111111111111111111111111111111101111111011111111111111101111111111011111110111111111111111111010111101111111111111110111111101111110111111110111111011011111111111111111111111111101111101111001111111111001111111111111111111111110011101111111111111110011111111111101111011111111001111110111111111111011110111111111111111111111111101111001111111111111111101111001011111111011111101111111011111010111111111111111110111111111111111111101111111101111111111111111111111011111111111011110111111111111111111111111111111111101;
    assign test_vec[91] = 1024'b1010111110111110111111111111111010011111111110111111111001111111111111111111110111111111111111011111111111011111111111111111111111111111111111111111111101111111111111111111111011110111111111101111111111111101111111111111111010011011000111111101111111011111111101111111111110111111111011111111111111101111111111111111111111111111101111111111111111111111111111111111111011111111111110111001111111110111111111111111111101011111111101111011111111011101111111111001111111111111111111111111111111100101111111011111111111010111111111110111111111111111111111111111111110111111111101111111111111111111111111111101110111111111111111111111111111111111111111111111011111101111111111111101111111111110111111111100111111111111101111010101111110110111111111111111111111111101101111111101110110110111111111111111111111111111111111111111111111111111111011111111011111111111110111111111111011111111110111111111111110011110110111111101111111111111111111111111111110100111111111111110111111011001111111111111111111111110111111111111111111111101;
    assign test_vec[92] = 1024'b0111111011111110101111111111101111111111111111111110111110011111111111111111110111111111111111010011111011111111100111101110110101011111111111011111111111111111111111110111111111111111111011101111111111111110011001111111111111111111111111111101111111110111101111111101111111101111111011110111111101111111111111111111111111011110111110111011111111111111111111111111111011111111111111101111111111111111111111111111111111101101111111111111110111111111111111111111111111111101001111111111111111111111111111111111111111111111111111110111011111111111110011111111111111111111111111111111111111111111111111111111111111111011111111111101111111111111111101111111111011111001111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111011110111010111111111111111111110111111111111111111011111111111111010111111111111101101011111111111011101111110111111111111111111011111011111111111110111111111111111111011111111111111111111111111111111111111111101111111111111111110111111111111111101111111101101111111;
    assign test_vec[93] = 1024'b1111111011111111111110111111011011011111111111111111111011111111101111111111111111111111111110111101111110111101011101111111111111101111101011111111111111111111011111111111111111110111111111111111111111111111111111111111111111111111101111110111111111111111111111111101111111111111111111111111111111101111111111111111111111111111011111111111110111111111111111111111111111111101001111111111111111111111111111001101111101111111111111111111101111111111111111111111111111101111101111111111111111111111111111111111111111011111111111111111111111111111111111111110111111111110101111111110101111111111111111111111111111111111111101011111111110111111001111111111111111111111101111111111111011110111111111110110111111011111100111111111111111111111111111111111111111111110111111111101111111111111111111111111111111111111011111111111111111111011111111111111111111111111111110111101111011011011111111111111111111111111111111111111111101111111111111010111111111111111011111110111101111111101111111111111101111111111111111111111101110111111;
    assign test_vec[94] = 1024'b1111111111111111111111111111111111111111111111111111101011111111010111111110111111111111111111111111111111111110111111011111111111111101111111111101101111111111111011111111111111111111111011111111111111111111111101111111111111111111011111111111111111111111111111111001111111111111101011111111111111011111011011111101111111011111111111101111111101111011111111111111111111111111101110111111111111111110111011101111111011111111101111111101111111111110111110111111111111111110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111110011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111101111111011111111110110111111111111111101111111111111111110111111111111111111111111111110111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111101011111110111111111110111111111111111111111111111111111111110111110111111111111111111111111111011111101111111111111111111101111110111111111;
    assign test_vec[95] = 1024'b1011111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111110011111111111111111111111111111111111111111111111111111111111111010111111111111111101111111111111111111011111111111111011111111111111111111110111111101101111111111111111111111111111111111111111111101011111011111101111111011111111111111111111111111100001111111110011111111111111100111111111111111111111110111111111111111111111111111011011111111101011111111111101011111111111011111111111111111111111111111111111011111111111111111011111111111111111111111111101011111111111111111111111111101111110111111111111011111110111111111111111101111111111111111111111111111111111111111111111111111111110111101111111111111101111111111111111111111111110111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111011111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111110111111011111111111;
    assign test_vec[96] = 1024'b1111101101111111111111111111111111111110111111111111111111101111111111111111111011111111111111111111111111110111111111111111111111111111111111111111101111111111111111111111111101011111111111111111111111111111110110111111111111111110111111111111111111111111011011011111111110111111011111111111111111111111111111111111101111111111111111111111111111111011111111111111111111111111111111101111111111111110111111111111101111011101111111101111111111111110111111111111111111111111111111111011111111111111111111111101111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111011111111011111111111111111111111111111111111101111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111110111111101111111111111111111111111111111111111111111111111111111111101111111111110111110111111111111111111;
    assign test_vec[97] = 1024'b1111111111111111111111110111111011111110111111111111111111110111111111110111111101111111111111111111111111111111110111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111111011111111011111111110101111111111111111111111111111111111111111111111110111111111111111110111111111111111111111111111111011111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111110111111111111111111101101111111111111111111111111111111111011111111011111111111111111111111111111111111111110111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111110111111111101111101;
    assign test_vec[98] = 1024'b1111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111011111011111111111111111111111111111111111111111110111110111111111111111111111111111111111111111111111111111101111111111111111111111111101111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111001110111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111101111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111;
    assign test_vec[99] = 1024'b1111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111110111111111111111111111111111111111111111101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111;
    assign test_vec[100] = 1024'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

    assign deque = full && !empty;
    assign debug_mode = '0;
    assign spi_reg_lsb = '0;

    logic [9:0] count, latch_count;
    logic [31:0][1023:0] temp0, temp1;
    logic [1023:0] temp2;

    always_ff @(posedge clk) begin
        // for (int i = 0; i < es_sources; i++) begin
        //     ES_in[i] <= $urandom_range(0,1);
        // end
        if (rst) begin
            for (int i = 0; i < es_sources; i++) begin
                ES_in[i] <= test_vec[100][0];  // this is your biased input and then adjust to calibration after
                temp0[i] <= '0;
                temp1[i] <= '0;
            end
            temp2 <= '0;
            count <= '0;
            latch_count <= '0;
            
        end else if (count == 1023) begin
            for(int i = 0; i < latch_sources; i++) begin
                // temp0[i] <= test_vec[arr_n[i]* 1.5625];
                // temp1[i] <= test_vec[arr_p[i]* 1.5625];
                int idx_n, idx_p;
                idx_n = int'(arr_n[i] * 1.5625);
                idx_p = int'(arr_p[i] * 1.5625);
                // temp0[i] <= test_vec[100 - idx_n];
                // temp1[i] <= test_vec[idx_p];
                // temp2 <= temp1 + temp0;
                temp2 <= (idx_p - idx_n < 0) ? '0 : (idx_p - idx_n) / 2;
                ES_in[i] <= test_vec[temp2][latch_count];
            end
            latch_count <= latch_count+1;

        end else begin
            count <= count + 1;
        end
    end

    oht_top dut (
        .clk(clk),
        .rst(rst),

        .ES_in(ES_in),
        .deque(deque),
        .debug_mode(debug_mode),
        .spi_reg_lsb(spi_reg_lsb),

        .cond_out(cond_out),
        .full(full),
        .empty(empty),
        .arr_n(arr_n),
        .arr_p(arr_p),
        .j_disable_arr(j_disable_arr),
        .rd_good_arr(rd_good_arr)

    );

    initial begin
		$fsdbDumpfile("oht_top_dump.fsdb");
		$fsdbDumpvars(0, "+all");
		rst = 1'b1;
        // if (rst) begin
        //     for (int i = 0; i < es_sources; i++) begin
        //         ES_in[i] = test_vec[100][0];  // this is your biased input and then adjust to calibration after
        //     end
        //     count = '0;
        //     latch_count = '0;
        // end

        #10ns
		rst = 1'b0;
        // forever begin
        //     #1ns;
        //         for(int i = 0; i < latch_sources; i++) begin
        //             ES_in[i] <= test_vec[arr_n[i]][latch_count];
        //         end
        //         latch_count <= latch_count+1;
        //         if (latch_count == 1023) break;
        //     #1ns;
        // end
		#100000ns
		$finish();
	end

endmodule

